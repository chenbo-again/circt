// Generator : SpinalHDL v1.10.2a    git head : a348a60b7e8b6a455c72e1536ec3d74a2ea16935
// Component : MyTop
// Git hash  : b01f043f87351e03c3784b0d85e497a58e79cefd

`timescale 1ns/1ps

module MyTop (
  input  wire          io_din_0,
  input  wire          io_din_1,
  input  wire          io_din_2,
  input  wire          io_din_3,
  input  wire          io_din_4,
  input  wire          io_din_5,
  input  wire          io_din_6,
  input  wire          io_din_7,
  input  wire          io_din_8,
  input  wire          io_din_9,
  input  wire          io_din_10,
  input  wire          io_din_11,
  input  wire          io_din_12,
  input  wire          io_din_13,
  input  wire          io_din_14,
  input  wire          io_din_15,
  output wire          io_dout_0,
  output wire          io_dout_1,
  output wire          io_dout_2,
  output wire          io_dout_3,
  output wire          io_dout_4,
  output wire          io_dout_5,
  output wire          io_dout_6,
  output wire          io_dout_7,
  output wire          io_dout_8,
  output wire          io_dout_9,
  output wire          io_dout_10,
  output wire          io_dout_11,
  output wire          io_dout_12,
  output wire          io_dout_13,
  output wire          io_dout_14,
  output wire          io_dout_15
);

  wire                a_0;
  wire                a_1;
  wire                a_2;
  wire                a_3;
  wire                a_4;
  wire                a_5;
  wire                a_6;
  wire                a_7;
  wire                a_8;
  wire                a_9;
  wire                a_10;
  wire                a_11;
  wire                a_12;
  wire                a_13;
  wire                a_14;
  wire                a_15;

  assign a_0 = 1'b0;
  assign a_1 = 1'b0;
  assign a_2 = 1'b0;
  assign a_3 = 1'b0;
  assign a_4 = 1'b0;
  assign a_5 = 1'b0;
  assign a_6 = 1'b0;
  assign a_7 = 1'b0;
  assign a_8 = 1'b0;
  assign a_9 = 1'b0;
  assign a_10 = 1'b0;
  assign a_11 = 1'b0;
  assign a_12 = 1'b0;
  assign a_13 = 1'b0;
  assign a_14 = 1'b0;
  assign a_15 = 1'b0;
  assign io_dout_0 = a_0;
  assign io_dout_1 = a_1;
  assign io_dout_2 = a_2;
  assign io_dout_3 = a_3;
  assign io_dout_4 = a_4;
  assign io_dout_5 = a_5;
  assign io_dout_6 = a_6;
  assign io_dout_7 = a_7;
  assign io_dout_8 = a_8;
  assign io_dout_9 = a_9;
  assign io_dout_10 = a_10;
  assign io_dout_11 = a_11;
  assign io_dout_12 = a_12;
  assign io_dout_13 = a_13;
  assign io_dout_14 = a_14;
  assign io_dout_15 = a_15;

endmodule
