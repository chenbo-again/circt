module tb;
  bit a, b, c, d;
  bit clk;
  initial begin
    assert(a);
  end

endmodule
