module string_ex ();

initial begin

end

endmodule